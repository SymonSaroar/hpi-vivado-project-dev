`timescale 1 ps / 1 ps

module design_wrapper
   (output_data_0);
  output [191:0]output_data_0;

  wire [191:0]output_data_0;

  design_1 design_1_i
       (.output_data_0(output_data_0));
endmodule
